--TYPE PACKAGE

package type_pkg is

	type lfo_shape_t is (SQUARE, TRI,SAW); 
	end package type_pkg;