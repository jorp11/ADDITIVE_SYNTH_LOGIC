-- clk_div_tb.vhd
